module clk_buffer(input mclk,output bclk);
buf d1 (bclk,mclk);

endmodule